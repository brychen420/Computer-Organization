module ALU_Ctrl( funct_i, ALUOp_i, ALU_operation_o, FURslt_o );

//I/O ports 
input      [6-1:0] funct_i;
input      [3-1:0] ALUOp_i;

output     [4-1:0] ALU_operation_o;  
output     [2-1:0] FURslt_o;
     
//Internal Signals
reg	    [4-1:0] ALU_operation_o;
wire	[2-1:0] FURslt_o;

//Main function
/*your code here*/

assign FURslt_o = ((funct_i == 6'b000000) || (funct_i == 6'b000010)) ? 2'b01 : 2'b00;
//Select exact operation
always@(*)begin
	if(ALUOp_i == 3'b010)begin
          case(funct_i)
            6'b010010: ALU_operation_o = 4'b0010; // add
			6'b010000: ALU_operation_o = 4'b0110; // sub
			6'b010100: ALU_operation_o = 4'b0001; // and
			6'b010110: ALU_operation_o = 4'b0000; // or
			6'b010101: ALU_operation_o = 4'b1100; // nor
			6'b100000: ALU_operation_o = 4'b0111; // slt
			6'b000000: ALU_operation_o = 4'b0001; // sll
			6'b000010: ALU_operation_o = 4'b0000; // srl
			default: ALU_operation_o = 4'b0000;
          endcase
        end
	else if(ALUOp_i == 3'b011)	ALU_operation_o = 4'b0010; //addi
	else if(ALUOp_i == 3'b001)	ALU_operation_o = 4'b0110; //beq (sub)
	else if(ALUOp_i == 3'b000)	ALU_operation_o = 4'b0010; //lw sw
	else if(ALUOp_i == 3'b110)	ALU_operation_o = 4'b1010; //bne
end

endmodule     
